module sign_extend(
    input  logic [31:0] instr,
    input  logic        ImmSrc,
    output logic [31:0] ImmOp
);



endmodule