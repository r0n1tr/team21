module top_pc #(
    parameter ADDRESS_WIDTH = 32,
              DATA_WIDTH = 32
)(
    input  logic                  clk,
    input  logic                  rst,
    input  logic                  trigger,
    input  logic [1:0]            pcsrc,
    input  logic [DATA_WIDTH-1:0] immext,
    input  logic [DATA_WIDTH-1:0] aluresult,
    
    output logic [ADDRESS_WIDTH-1:0] pcplus4,  // output this for use in result_mux (for jal instruction)
    output logic [ADDRESS_WIDTH-1:0] pctarget, // output this for use in result_mux (for auipc instruction)
    output logic [ADDRESS_WIDTH-1:0] pc
);

logic [ADDRESS_WIDTH-1:0] next_pc;

pc_reg pc_reg(
    .clk(clk),
    .next_pc(next_pc),
    
    .pc(pc)
);

pc_mux pc_mux (
    .aluresult(aluresult),
    .immext(immext),
    .pc(pc),
    .pcsrc(pcsrc),
    .rst(rst),
    .trigger(trigger),
    
    .pcplus4(pcplus4),
    .pctarget(pctarget),
    .next_pc(next_pc)
);

endmodule
