module topalu #(
    
) (
    input logic AD1,
    input logic AD2,
    input logic AD3,
    input logic WE3,
    input logic WD3,
    input logic clk,
    output logic EQ,
    output logic ALUout
);

regfile myregfile(

)

mux mymux(

)

alu myalu(

)
    
endmodule